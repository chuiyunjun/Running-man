module datapath(input clk,	reset_n, drawing_floors, draw_man, erase, x_original, y_original, normal1crouch0,
						output reg draw_floors_finish,
						output reg draw_man_finish,
						output reg erase_finish,
						output reg [2:0] color,
						output reg [7:0] x,
						output reg [6:0] y);
				
				
				
						
				always @(posedge clk)
				begin
					if(!reset_n)
						begin
							x <= 8'd0;
							y <= 7'd35;
						end
					else if(drawing_floors)
						begin
							color = 3'b101;
							if(x == 8'd159)
								begin
									x <= 0;
									if(y >= 7'd35 && y <= 7'd38 || y >= 7'd75 && y <= 7'd78 || y >= 7'd115 && y <= 7'd118)
										begin y <= y + 1; end 
									else if (y == 7'd39 || y == 7'd79)
										begin y <= y + 40; end
									else if (y == 7'd119)
										begin draw_floors_finish <= 1; end
								end
							else
								begin
									x <= x + 1;
								end
						end
					else if(draw_man || erase)
						color = draw_man ? 3'b111:3'b000;
						begin
							begin
									if(q == 6'd0) begin
										x = x_original + 2'd3;
										y = y_original;
									end	
									else if (q == 6'd1) begin
										x = x_original + 3'd4;
										y = y_original;
									end
									else if(q == 6'd2) begin
										x = x_original + 3'd5;
										y = y_original;
									end
									else if(q == 6'd3) begin
										x = x_original + 2'd3;
										y = y_original + 1'b1;
									end	
									else if(q == 6'd4) begin
										x = x_original + 3'd5;
										y = y_original + 1'd1;
									end
									else if(q == 6'd5) begin
										x = x_original + 2'd3;
										y = y_original + 2'd2;
									end	
									else if(q == 6'd6) begin
										x = x_original + 3'd4;
										y = y_original + 2'd2;
									end	
									else if(q == 6'd7) begin
										x = x_original + 3'd5;
										y = y_original + 2'd2;
									end
									else if(q == 6'd8) begin
										x = x_original;
										y = y_original + 3'd3;
									end
									else if(q == 6'd9) begin
										x = x_original + 1'd1;
										y = y_original + 3'd3;
									end
									else if(q == 6'd10) begin
										x = x_original + 2'd2;
										y = y_original + 3'd3;
									end
									else if(q == 6'd11) begin
										x = x_original + 2'd3;
										y = y_original + 3'd3;
									end
									else if(q == 6'd12) begin
										x = x_original;
										y = y_original + 3'd4;
									end
									else if(q == 6'd13) begin
										x = x_original + 1'd1;
										y = y_original + 3'd4;
									end
									else if(q == 6'd14) begin
										x = x_original + 2'd2;
										y = y_original + 3'd4;
									end
									else if(q == 6'd15) begin
										x = x_original + 2'd3;
										y = y_original + 3'd4;
									end	
									else if(q == 6'd16) begin
										x = x_original;
										y = y_original + 3'd5;
									end
									else if(q == 6'd17) begin
										x = x_original + 1'd1;
										y = y_original + 3'd5;
									end
									else if(q == 6'd18) begin
										x = x_original + 2'd2;
										y = y_original + 3'd5;
									end
									else if(q == 6'd19) begin
										x = x_original + 3'd3;
										y = y_original + 3'd5;
									end
									else if(q == 6'd20) begin
										x = x_original;
										y = y_original + 3'd6;
									end	
									else if(q == 6'd21) begin
										x = x_original + 3'd3;
										y = y_original + 3'd6;
									end
									else if(q == 6'd22) begin
										x = x_original - 1'd1;
										y = y_original + 2'd3;
									end
									else if(q == 6'd23) begin
										x = x_original - 2'd2;
										y = y_original + 2'd3;
									end
									else if(q == 6'd24) begin
										x = x_original + 2'd3;
										y = y_original - 1'd1;
									end
									else if(q == 6'd25) begin
										x = x_original + 3'd5;
										y = y_original - 1'd1;

									end

								end
						end
				end
				
				reg [5:0] q;
				always @(clk)
				begin
					if(!resetn)
						begin
							draw_man_finish <= 0;
							erase_finish <= 0;
							q <= 0;
						end

					if(q == 6'd25)
						begin
							q <= 0;
							if(draw_man)
								begin
									draw_man_finish <= 1;
									erase_finish <= 0;
									draw_floors_finish <= 0;
								end
							else if(erase)
								begin
									erase_finish <= 1;
									draw_man_finish <= 0;
								end
						end
					else
						begin
							q <= q + 1;
						end
				end
						
endmodule